*** SPICE deck for cell inv_1211753{lay} from library inverter_1211753
*** Created on Sun Dec 14, 2025 18:33:03
*** Last revised on Mon Dec 15, 2025 19:49:59
*** Written on Mon Dec 15, 2025 20:13:29 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: inverter_1211753:inv_1211753{lay}
Mnmos_1 0 A Y 0 NMOS L=0.4U W=2U AS=7.68P AD=11.08P PS=20U PD=24.8U
Mpmos_1 vdd A Y vdd PMOS L=0.4U W=6U AS=7.68P AD=29.48P PS=20U PD=56.8U

* Spice Code nodes in cell cell 'inverter_1211753:inv_1211753{lay}'
VDD  vdd 0 DC 5
VIN  A   0 PWL(10n 0  20n 5  50n 5  60n 0)
CLOAD Y  0 250f
; Fall time of V(Y): 90% -> 10% (4.5V to 0.5V) around the first transition
.measure tran tf  TRIG v(Y) VAL=4.5 FALL=1 TD=8n  TARG v(Y) VAL=0.5 FALL=1
; Rise time of V(Y): 10% -> 90% (0.5V to 4.5V) around the second transition
.measure tran tr  TRIG v(Y) VAL=0.5 RISE=1 TD=50n TARG v(Y) VAL=4.5 RISE=1
; (optional but recommended) propagation delays at 50% VDD (2.5V)
.measure tran tphl TRIG v(A) VAL=2.5 RISE=1          TARG v(Y) VAL=2.5 FALL=1
.measure tran tplh TRIG v(A) VAL=2.5 FALL=1          TARG v(Y) VAL=2.5 RISE=1
.tran 0 0.1u
.include "C:\ltspice\C5_models.txt"
.END
