*** SPICE deck for cell triple_and{sch} from library application
*** Created on Mon Dec 15, 2025 18:15:05
*** Last revised on Tue Dec 16, 2025 02:50:45
*** Written on Tue Dec 16, 2025 03:02:17 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT inverter_1211753__inv_1211753 FROM CELL inverter_1211753:inv_1211753{sch}
.SUBCKT inverter_1211753__inv_1211753 A Y
** GLOBAL 0
** GLOBAL vdd
Mnmos_0 Y A 0 0 NMOS L=0.4U W=2U
Mpmos_0 vdd A Y vdd PMOS L=0.4U W=6U
.ENDS inverter_1211753__inv_1211753

*** SUBCIRCUIT nand_2_1211753__nand_1211753 FROM CELL nand_2_1211753:nand_1211753{sch}
.SUBCKT nand_2_1211753__nand_1211753 A B Y
** GLOBAL 0
** GLOBAL vdd
Mnmos_0 net_0 B 0 0 NMOS L=0.4U W=4U
Mnmos_1 Y A net_0 0 NMOS L=0.4U W=4U
Mpmos_0 vdd A Y vdd PMOS L=0.4U W=6U
Mpmos_1 vdd B Y vdd PMOS L=0.4U W=6U
.ENDS nand_2_1211753__nand_1211753

*** SUBCIRCUIT NOR_3_1211753__nor_1211753 FROM CELL NOR_3_1211753:nor_1211753{sch}
.SUBCKT NOR_3_1211753__nor_1211753 A B C Y
** GLOBAL 0
** GLOBAL vdd
Mnmos_0 Y A 0 0 NMOS L=0.4U W=2U
Mnmos_1 Y B 0 0 NMOS L=0.4U W=2U
Mnmos_2 Y C 0 0 NMOS L=0.4U W=2U
Mpmos_0 net_13 A Y vdd PMOS L=0.4U W=18U
Mpmos_1 net_14 B net_13 vdd PMOS L=0.4U W=18U
Mpmos_2 vdd C net_14 vdd PMOS L=0.4U W=18U
.ENDS NOR_3_1211753__nor_1211753

.global 0 vdd

*** TOP LEVEL CELL: triple_and{sch}
Xinv_1211_0 C net_10 inverter_1211753__inv_1211753
Xnand_121_0 A B net_12 nand_2_1211753__nand_1211753
Xnor_1211_0 net_12 net_10 0 Y NOR_3_1211753__nor_1211753

* Spice Code nodes in cell cell 'triple_and{sch}'
VDD  vdd 0 DC 5
VA  A 0 PWL(10n 0  20n 5  50n 5  60n 0)
VB  B 0 PWL(15n 0  25n 5  55n 5  65n 0)
VC  C 0 PWL(30n 0  40n 5  70n 5  80n 0)
CLOAD Y  0 250ff
.measure tran tf  TRIG v(Y) VAL=4.5 FALL=1 TD=8n  TARG v(Y) VAL=0.5 FALL=1
.measure tran tr  TRIG v(Y) VAL=0.5 RISE=1 TD=50n TARG v(Y) VAL=4.5 RISE=1
.measure tran tphl TRIG v(A) VAL=2.5 RISE=1          TARG v(Y) VAL=2.5 FALL=1
.measure tran tplh TRIG v(A) VAL=2.5 FALL=1          TARG v(Y) VAL=2.5 RISE=1
.tran 0.1u
.include "C:\ltspice\C5_models.txt"
.END
