*** SPICE deck for cell inv_1211753{sch} from library inverter_1211753
*** Created on Sun Dec 14, 2025 16:22:37
*** Last revised on Tue Dec 16, 2025 02:48:24
*** Written on Tue Dec 16, 2025 02:48:33 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global 0 vdd

*** TOP LEVEL CELL: inverter_1211753:inv_1211753{sch}
Mnmos_0 Y A 0 0 NMOS L=0.4U W=2U
Mpmos_0 vdd A Y vdd PMOS L=0.4U W=6U

* Spice Code nodes in cell cell 'inverter_1211753:inv_1211753{sch}'
VDD  vdd 0 DC 5
VIN  A   0 PWL(10n 0  20n 5  50n 5  60n 0)
CLOAD Y  0 250ff
.measure tran tf  TRIG v(Y) VAL=4.5 FALL=1 TD=8n  TARG v(Y) VAL=0.5 FALL=1
.measure tran tr  TRIG v(Y) VAL=0.5 RISE=1 TD=50n TARG v(Y) VAL=4.5 RISE=1
.measure tran tphl TRIG v(A) VAL=2.5 RISE=1          TARG v(Y) VAL=2.5 FALL=1
.measure tran tplh TRIG v(A) VAL=2.5 FALL=1          TARG v(Y) VAL=2.5 RISE=1
.tran 0 0.1u
.include "C:\ltspice\C5_models.txt"
.END
